module main

import naml

fn main() {
	println(naml.read_file('./test.naml') ? )
}